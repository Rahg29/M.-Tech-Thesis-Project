`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 10.09.2018 18:58:56
// Design Name: 
// Module Name: AIM
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module dim8(
input signed [8:0] A1, A2, A3, A4, A5, A6, A7, A8,
input signed [1:0] W1, W2, W3, W4, W5, W6, W7, W8,
input clk,
output reg signed [11:0] out_neuron
);

reg [7:0] Act_Index;
reg [7:0] Weight_Index;

reg signed [8:0] Activation [0:7];
reg signed [1:0] Weight [0:7];

reg [4:0] Inc_Act [0:7];
reg [4:0] Inc_Weight [0:7];

reg signed [8:0] Act_element [0:5];
reg signed [8:0] Weight_element [0:5];

reg [7:0] and_op;

integer i= 0, c= 0, f= 0, e= 0, g= 0, reset = 1;

reg signed [11:0] y= 12'd0;

reg [1:0]Pres_state;
reg [1:0] Next_state;

parameter S0=2'd0;
parameter S1=2'd1;
parameter S2=2'd2;
parameter S3=2'd3;

always @(posedge clk)
begin
    if (reset == 1'd1)
    Pres_state = S0;
    
    else
    Pres_state = Next_state;
end


always @(posedge clk)
begin

case(Pres_state)

S0:begin
reset=0;

Weight[0] = W1;
Weight[1] = W2;
Weight[2] = W3;
Weight[3] = W4;
Weight[4] = W5;
Weight[5] = W6;
Weight[6] = W7;
Weight[7] = W8;

Activation[0] = A1;
Activation[1] = A2;
Activation[2] = A3;
Activation[3] = A4;
Activation[4] = A5;
Activation[5] = A6;
Activation[6] = A7;
Activation[7] = A8;

Next_state = S1;
end


S1:begin
    //reset=1'd0;
    out_neuron[11:0] = i;
    if (i<=7)
    begin
     
        if(Weight[i] == 2'd0 && Activation[i] == 9'd0)
            begin
            Weight_Index[i] = 1'b0;
            Act_Index[i] = 1'b0;
            c = c + Act_Index[i];
            f = f + Weight_Index[i];
            Inc_Act[i] = c;
            Inc_Weight[i] = f;
            i = i+1;
            Next_state = S1;
            end
            
            else if(Weight[i] == 2'd0)
            begin
            Weight_Index[i] = 1'b0;
            Act_element[e] = Activation[i];
            Act_Index[i] = 1'b1;
            c = c + Act_Index[i];
            f = f + Weight_Index[i];
            Inc_Act[i] = c;
            Inc_Weight[i] = f;
            i = i+1;
            e = e+1;
            Next_state = S1;
            end
            
            else if(Activation[i] == 9'd0)
            begin
            Act_Index[i] = 1'b0;
            Weight_Index[i] = 1'b1;
            Weight_element[g] = Weight[i];
            c = c + Act_Index[i];
            f = f + Weight_Index[i];
            Inc_Act[i] = c;
            Inc_Weight[i] = f;
            g = g+1;
            i = i+1;
            Next_state = S1;
            end
            
            else
            begin
            Act_element[e] = Activation[i];
            Weight_element[g] = Weight[i];
            Act_Index[i] = 1'b1;
            Weight_Index[i] = 1'b1;
            c = c + Act_Index[i];
            f = f + Weight_Index[i];
            Inc_Act[i] = c;
            Inc_Weight[i] = f;
            i = i+1;
            e = e+1;
            g = g+1;
            Next_state = S1;
            end         
    end
    
    else 
    begin
    Next_state = S2;
    end
end


S2: begin
    and_op = Act_Index & Weight_Index;
    out_neuron[11:0] = 12'd10;
    i=0;
    Next_state = S3;
    end

S3:begin
    out_neuron[11:0] = 20 + i;
    if (i<=7)
        begin
            if(and_op[i] == 1'b1)
            begin
            y = y + Weight_element[Inc_Weight[i]-1] * Act_element[Inc_Act[i]-1];
            i = i+1;
            Next_state = S3;
            end
            
            else
            begin
            i = i+1;
            Next_state = S3;
            end
        end
        
    else
    out_neuron[11:0] = y[11:0];
  end


endcase
end


endmodule
